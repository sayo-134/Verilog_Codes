module stimulus;

reg clk;
reg reset;  
wire[3:0] q;  
  
  
  
